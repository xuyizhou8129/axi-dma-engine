// optional skid buffer / small FIFO

