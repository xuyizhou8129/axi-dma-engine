// optional 64↔32 packing/unpacking

