// top wrapper: AXI-Lite slave + DMA engine + IRQ

