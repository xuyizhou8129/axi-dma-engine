// FIFO: decoupling buffers for descriptor queue, read data, writeback

