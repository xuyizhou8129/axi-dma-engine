// Descriptor fetch: AXI4 read to pull descriptors from system memory

