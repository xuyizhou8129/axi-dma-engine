// SRAM controller: converts stream data into SRAM write/read cycles, handles timing/masking

