// simple AXI memory model

