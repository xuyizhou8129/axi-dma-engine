// AXI4 read address/data channel handling

