// optional (if multi-channel)

