// reg decode + fields + reset values

