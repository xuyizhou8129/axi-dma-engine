// high-level FSM: IDLE→READ→WRITE→DONE

