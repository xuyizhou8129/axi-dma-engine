// done/error pending/mask + irq output

