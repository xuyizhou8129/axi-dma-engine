// AXI4 write address/data/resp handling

