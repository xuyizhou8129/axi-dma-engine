// Scheduler / Control FSM: pops descriptors, validates, orchestrates transaction sequence

