// typedefs/params (desc format, enums)

