// Descriptor queue/FIFO: buffers fetched descriptors for scheduler

