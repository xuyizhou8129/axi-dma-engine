// Ring manager: tracks head/tail, computes descriptor addresses, handles wraparound

