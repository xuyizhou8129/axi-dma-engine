// Data mover: coordinates AXI read/write engines and SRAM controller for payload transfer

