// SRAM signals + adapter

