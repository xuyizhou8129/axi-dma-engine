// AXI4-Lite register bank

