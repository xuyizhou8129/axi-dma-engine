// AXI4-Lite register bank + reg decode + fields + reset values

